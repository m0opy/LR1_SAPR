module apb_slave

(
  input pclk, 			// ????????????
  input presetn, 		// ?????? ?????? (?????????)
  input [31:0] paddr, 		// ????? ?????????
  input [31:0] pwdata, 		// ?????? ??? ??????
  input psel, 			// ??????? ?????? ?????????
  input penable, 		// ??????? ???????? ??????????
  input pwrite, 		// ??????? ???????? ??????
  output logic pready, 		// ??????? ?????????? ?? ??????????
  output logic pslverr, 	// ???????????? ??????: ??????? ?????? ??? ?????????
  output logic [31:0] prdata 	// ??????????? ??????
);

logic [31:0] reg_group;   	// 0x00
logic [31:0] reg_date;          // 0x04
logic [31:0] reg_surname;       // 0x08
logic [31:0] reg_name;          // 0x0C

//APB FSM
enum logic [1:0] {
  APB_SETUP,	// ???? ??????????
  APB_W_ENABLE,	// ???? ??????
  APB_R_ENABLE	// ???? ??????
} apb_st;

always @(posedge pclk)		// ???????????? ?? ????? ?????
  if (!presetn)			// ???? ?????? ?????? -- ???????? ???????? ????????? ????????
  begin
    // ????????? ?????????
    prdata <= '0;			
    pslverr <= 1'b0;		
    pready <= 1'b0;			
    reg_group <= 32'h0;
    reg_date <= 32'h0;
    reg_surname <= 32'h0;
    reg_name <= 32'h0;
    apb_st <= APB_SETUP;	// ????????? ??????????
  end
  else				// ???? ?? ?????
  begin
    case(apb_st)
      APB_SETUP:		// ????????? ??????????
      begin: apb_setup_st
	prdata <= '0;		// ????? ??????
	pslverr <= 1'b0;	// ????? ??????
	pready <= 1'b0;		// ?????????? ?? ??????
	// ENABLE => PSEL = 1(?????????? ??????) && PENABLE = 0(?????????? ?? ???????)
	if (psel && !penable)
	begin
	  if (pwrite == 1'b1)	    // ???????? ??????
	  begin
	    apb_st <= APB_W_ENABLE; // ??????? ? ???? ??????
	  end
	else			    // ???????? ??????
	begin
	  apb_st <= APB_R_ENABLE;   // ??????? ? ???? ??????
	end
      end
    end: apb_setup_st

  // ???? ??????
  APB_W_ENABLE:
  begin: apb_w_en_st
    // ???? ?????????? ??????, ??????? ?????????? ? ???????? ??????
    if (psel && penable && pwrite)
    begin
      pready <= 1'b1; // ?????????? ??????????
      case (paddr[7:0])
        8'h0: begin
	  // ?????? ? ??????? ?? ????????? 0
	  reg_group <= pwdata;
	  $display("[%0t] APB WRITE  0x00 <= 0x%08h (GROUP)",   $time, pwdata);
	end

	8'h4: begin
	  // ?????? ? ??????? ?? ????????? 4
	  reg_date <= pwdata;
	  $display("[%0t] APB WRITE  0x04 <= 0x%08h (DATE)", $time, pwdata);
	end

	8'h8: begin
	  // ?????? ? ??????? ?? ????????? 8
	  reg_surname <= pwdata;
	  $display("[%0t] APB WRITE  0x08 <= 0x%08h (SUR)", $time, pwdata);
	end

	8'h0C: begin
	  // ?????? ? ??????? ?? ????????? 12
	  reg_name <= pwdata;
	  $display("[%0t] APB WRITE  0x0C <= 0x%08h (NAME)",$time, pwdata);
	end

	default:
	begin
	  // ???? ??????
	  pslverr <= 1'b1;
	  $display("[%0t] APB WRITE  ERROR bad addr=0x%08h", $time, paddr);
	end
      endcase
      apb_st <= APB_SETUP; // ??????????? ? ???????? ?????????
    end
  end: apb_w_en_st
  
  // ???? ??????
  APB_R_ENABLE:
  begin: apb_r_en_st
    // ???? ?????????? ??????, ??????? ?????????? ? ???????? ??????
    if (psel && penable && !pwrite)
    begin
      pready <= 1'b1; // ?????????? ?????????? 
      case (paddr[7:0])
	8'h0: begin
	  // ?????? ?? ???????? ?? ????????? 0
	  prdata <= reg_group;
	  $display("[%0t] APB READ   0x00 => 0x%08h (GROUP)", $time, reg_group);
	end

	8'h4: begin
	  // ?????? ?? ???????? ?? ????????? 4
	  prdata <= reg_date;
	  $display("[%0t] APB READ   0x04 => 0x%08h (DATE)", $time, reg_date);
	end

	8'h8: begin
	  // ?????? ?? ???????? ?? ????????? 8
	  prdata <= reg_surname;
	  $display("[%0t] APB READ   0x08 => 0x%08h (SUR)",  $time, reg_surname);
 	end

	8'h0C: begin
	  // ?????? ?? ???????? ?? ????????? 12
	  prdata <= reg_name;
	  $display("[%0t] APB READ   0x0C => 0x%08h (NAME)", $time, reg_name);
 	end

	default:
	begin
	  pslverr <= 1'b1; // ???? ??????
	  $display("[%0t] APB READ   ERROR bad addr=0x%08h", $time, paddr);
	end
      endcase
      apb_st <= APB_SETUP; // ??????? ? ???????? ?????????
    end
  end: apb_r_en_st

  default:
  begin
    pslverr <= 1'b1; // ???? ??????
  end
endcase

end // ?????????? ???? ?????? always

endmodule



