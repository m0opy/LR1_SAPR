module TB;

logic pclk;		// ????????????
logic presetn;		// ?????? ?????? (?????????)
logic psel;		// ??????? ?????? ?????????
logic penable;		// ??????? ???????? ??????????
logic pwrite;		// ??????? ???????? ??????
logic [31:0] paddr;	// ????? ?????????
logic [31:0] pwdata;	// ?????? ??? ??????
wire [31:0] prdata;	// ??????????? ??????
wire pready;		// ??????? ?????????? ?? ??????????
wire pslverr;		// ???????????? ??????: ??????? ?????? ??? ?????????

parameter p_device_offset = 32'h7000_0000; // ??????? ????? ?????????? ? ???????? ????????????

logic [31:0] data_from_device; // ??????, ????????? ? ????

apb_slave DUT
(
  .pclk(pclk), 		// ??????????? ????? 		
  .presetn, 		// ????? (??????????? ?????? .presetn(presetn)) 		
  .paddr(paddr), 	// ????? 	
  .pwdata(pwdata), 	// ?????? ?? ??????	
  .psel(psel), 		// ????? ?????????? 		
  .penable(penable), 	// ???? ENABLE 	
  .pwrite(pwrite), 	// ???????? ??????/?????? 	
  .pready(pready), 	// ?????????? ??????????	
  .pslverr(pslverr), 	// ??????	
  .prdata(prdata) 	// ?????? ?? ??????	
);

localparam [31:0] A_GROUP = p_device_offset + 32'h00; 	// ???????? 0x00: ??????? �????? ? ??????�
localparam [31:0] A_DATE = p_device_offset + 32'h04; 	// ???????? 0x04: ??????? �????�
localparam [31:0] A_SUR = p_device_offset + 32'h08; 	// ???????? 0x08: ??????? �??????? (4 ASCII)�
localparam [31:0] A_NAME = p_device_offset + 32'h0C; 	// ???????? 0x0C: ??????? �??? (4 ASCII)�

localparam [31:0] STUDENT_GROUP = 32'd24; 	// ????? ? ??????
localparam [31:0] DATE = 32'h27102025; 		// ???? 
localparam [31:0] SUR  = {"S","H","C","H"}; 	// ?????? 4 ????? ??????? ? ASCII
localparam [31:0] NAME = {"P","O","L","I"}; 	// ?????? 4 ????? ????? ? ASCII

task apb_write(input [31:0] addr, input [31:0] data); // ?????????? ?????? ?? APB
  wait ((penable==0) && (pready == 0)); // ???????? ???????????? ????(penable==0) ? ??????????(pready == 0)
  @(posedge pclk); 		// ????
  psel <= 1'b1; 		// ????? ??????????
  paddr[31:0] <= addr[31:0]; 	// ?????????? ?????
  pwdata[31:0] <= data[31:0]; 	// ?????????? ?????? ?? ??????
  pwrite <= 1'b1; 		// ???????? ??????
 
  @(posedge pclk);		// ????
  penable <= 1'b1;		// ?????????? ??????????

  @(posedge pclk);		// ????
  wait (pready == 1'b1);	// ???? ?????????? ??????????

  @(posedge pclk);		// ????
  psel <= 1'b0;			// ??????????? ??????????
  penable <= 1'b0;		// ?????????? ?????????????
  pwrite <= 1'b0;		// ????????? ????????

  @(posedge pclk);		// ????
endtask


task apb_read(input [31:0] addr, output logic [31:0] data); // ?????????? ?????? ?? APB
  wait ((penable==0) && (pready == 0)); // ???????? ???????????? ????(penable==0) ? ??????????(pready == 0)

  @(posedge pclk); 		// ????
  psel <= 1'b1; 		// ????? ??????????
  pwrite <= 1'b0; 		// ???????? ??????
  paddr[31:0] <= addr[31:0]; 	// ??????????? ??????

  @(posedge pclk);		// ????
  penable <= 1'b1;		// ?????????? ??????????

  @(posedge pclk);		// ????
  wait (pready == 1'b1);	// ???? ?????????? ??????????
  data[31:0] = prdata[31:0];	// ?????? ??????

  @(posedge pclk);		// ????
  psel <= 1'b0;			// ???????????? ??????????
  penable <= 1'b0;		// ????? ??????????

  @(posedge pclk);		// ????
endtask

always
#10ns pclk=~pclk;  		// ????????? ????????? ???????

initial
begin
  // ?????????????
  pclk=0;
  presetn=1'b1; 
  psel='0; 
  penable='0;
  pwrite='0;
  paddr='0;
  pwdata='0;

  repeat (5) @(posedge pclk); 	// 5 ?????? ?? ??????
  presetn=1'b0; 		// ?????
  repeat (5) @(posedge pclk); 	// ????? 5 ??????
  presetn=1'b1; 		// ??????? ?????
  repeat (5) @(posedge pclk); 	// ?????? 5 ??????

  // ??????/?????? ?????? ?????? ? ??????
  apb_write(A_GROUP, STUDENT_GROUP);
  apb_read (A_GROUP, data_from_device);
  $display("GROUP wrote %0d, read %0d", STUDENT_GROUP, data_from_device);

  // ??????/?????? ???? ? ??????
  apb_write(A_DATE, DATE);
  apb_read (A_DATE, data_from_device);
  $display("DATE  wrote 0x%08h, read 0x%08h", DATE, data_from_device);

  // ??????/?????? 4-? ???? ??????? ? ??????
  apb_write(A_SUR, SUR);
  apb_read (A_SUR, data_from_device);
  $display("SUR   wrote 0x%08h, read 0x%08h", SUR, data_from_device);

  // ??????/?????? 4-? ???? ????? ? ??????
  apb_write(A_NAME, NAME);
  apb_read (A_NAME, data_from_device);
  $display("NAME  wrote 0x%08h, read 0x%08h", NAME, data_from_device);

  repeat (10) @(posedge pclk); // ????? ????? ????????
  $stop();
end

initial // ?????? ???????: ?????????? ????
begin   // ???????? ???????? ??? ?? ?????????
  $monitor("APB IF state: PENABLE=%b PREADY=%b PADDR=0x%h PWDATA=0x%h PRDATA=0x%h", penable, pready, paddr, pwdata, prdata);
end

endmodule // ????? ??????
