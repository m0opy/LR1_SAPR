module apb_slave

(
  input pclk, 			// ????????????
  input presetn, 		// ?????? ?????? (?????????)
  input [31:0] paddr, 		// ????? ?????????
  input [31:0] pwdata, 		// ?????? ??? ??????
  input psel, 			// ??????? ?????? ?????????
  input penable, 		// ??????? ???????? ??????????
  input pwrite, 		// ??????? ???????? ??????
  output logic pready, 		// ??????? ?????????? ?? ??????????
  output logic pslverr, 	// ???????????? ??????: ??????? ?????? ??? ?????????
  output logic [31:0] prdata 	// ??????????? ??????
);

logic [31:0] register_with_some_name;

//APB FSM
enum logic [1:0] {
  APB_SETUP,
  APB_W_ENABLE,
  APB_R_ENABLE
} apb_st;

always @(posedge pclk)		// ???????????? ?? ????? ?????
  if (!presetn)			// ???? ?????? ?????? -- ???????? ???????? ????????? ????????
  begin
    prdata <= '0;			
    pslverr <= 1'b0;		
    pready <= 1'b0;			
    register_with_some_name <= 32'h0;
    apb_st <= APB_SETUP;	// ????????? ??????????
  end
  else
  begin
    case(apb_st)
      APB_SETUP:
      begin: apb_setup_st
        // ???????? prdata ? pready (?????? ??????????)
	prdata <= '0;
	pready <= 1'b0;	
	// ENABLE => PSEL = 1 && PENABLE = 0
	if (psel && !penable)
	begin
	  if (pwrite == 1'b1)
	  begin
	    apb_st <= APB_W_ENABLE;
	  end
	else
	begin
	  apb_st <= APB_R_ENABLE;
	end
      end
    end: apb_setup_st

  APB_W_ENABLE:
  begin: apb_w_en_st
    // ??????????? ?????? ? ??????
    if (psel && penable && pwrite)
    begin
      pready <= 1'b1;
      case (paddr[7:0])
        8'h0: begin
	  // ?????? ? ??????? ?? ????????? 0
	  register_with_some_name <= pwdata;
	end

	8'h4: begin
	  // ?????? ? ??????? ?? ????????? 4
	end

	8'h8: begin
	  // ?????? ? ??????? ?? ????????? 8
	end

	default:
	begin
	  pslverr <= 1'b1;
	end
      endcase
      apb_st <= APB_SETUP;
    end
  end: apb_w_en_st

  APB_R_ENABLE:
  begin: apb_r_en_st
    if (psel && penable && !pwrite)
    begin
      pready <= 1'b1;
      case (paddr[7:0])
	8'h0: begin
	  // ?????? ?? ???????? ?? ????????? 0
	  prdata[31:0] <= register_with_some_name[31:0];
	end

	8'h4: begin
	  // ?????? ?? ???????? ?? ????????? 4
	end

	8'h8: begin
	  // ?????? ?? ???????? ?? ????????? 8
 	end

	default:
	begin
	  pslverr <= 1'b1;
	end
      endcase
      apb_st <= APB_SETUP;
    end
  end: apb_r_en_st

  default:
  begin
    pslverr <= 1'b1;
  end
endcase


// ????? ????????? ?????-?? ???????? ?????
//if (penable==1'b0)

if (register_with_some_name[0] == 1'b0)
begin
register_with_some_name <= 32'hAAAA_AAAA;
end
else
begin
register_with_some_name <= 32'h5555_5555;
end

end // ?????????? ???? ?????? always

endmodule



